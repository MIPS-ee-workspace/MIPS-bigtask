`timescale 1ns/1ns
module ALU_tb;

reg[31:0] _A;
reg[31:0] _B;
reg[5:0] _ALUFun;
reg _Sign;
wire[31:0] _Z;


ALU alu(.A(_A),.B(_B),.Sign(_Sign),.ALUFun(_ALUFun),.Z(_Z));

initial begin
	_Sign=1'b1;
	_ALUFun=6'd0;
	_A=32'b1000_0000_0000_0000_0000_0000_0000_0001;
	_B=32'b1000_0000_0000_0000_0000_0000_0000_0001;
	#100
	_Sign=1'b0;
	#100
	_Sign=1'b1;
	_ALUFun=1'b1;
	#100
	_A=32'b1000_0000_0000_0000_0000_0000_0000_0101;
	_B=32'b1000_0000_0000_0000_0000_0000_0000_0011;
	_ALUFun=6'b011000;
	#100
	_ALUFun=6'b011110;
	#100
	_ALUFun=6'b100000;
	_A[4:0]=5'b00100;
	_B=32'b1111_1111_1111_1111_1111_1111_1111_1111;
	#100
	_ALUFun=6'b100011;
	_A[4:0]=5'b00100;
	_B=32'b0111_1111_1111_1111_1111_1111_1111_1111;
	#100
	_ALUFun=6'b110011;
	_A=32'b1000_0000_0000_0000_0000_0000_0000_0001;
	_B=32'b1000_0000_0000_0000_0000_0000_0000_0001;
	#100
	_ALUFun=6'b111101;
	_A=32'b1000_0000_0000_0000_0000_0000_0000_0001;
	_B=32'b0000_0000_0000_0000_0000_0000_0000_0010;
	#100
	_ALUFun=6'b100011;
	_A[4:0]=5'b00100;
	_B=32'b1111_1111_1111_1111_1111_1111_1111_1111;
end


endmodule