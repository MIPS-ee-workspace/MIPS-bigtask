`timescale 1ns/1ps

module ROM (addr,data,overflow);
input [30:0] addr;
output [31:0] data;
output overflow;

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [31:0] ROM_DATA[ROM_SIZE-1:0];

assign data=(addr[30:2] < ROM_SIZE)?ROM_DATA[addr[30:2]]:32'b0;
assign overflow=(addr[30:2] >= ROM_SIZE)?1:0;

integer i;
initial begin

ROM_DATA[0] = 32'h08000003;
ROM_DATA[1] = 32'h0800000c;
ROM_DATA[2] = 32'h0800004f;
ROM_DATA[3] = 32'h3c104000;
ROM_DATA[4] = 32'h2008fff6;
ROM_DATA[5] = 32'hae080000;
ROM_DATA[6] = 32'hae080004;
ROM_DATA[7] = 32'h20080003;
ROM_DATA[8] = 32'hae080008;
ROM_DATA[9] = 32'h2004007c;
ROM_DATA[10] = 32'h200500a3;
ROM_DATA[11] = 32'h0800000b;
ROM_DATA[12] = 32'hafa10000;
ROM_DATA[13] = 32'hafa20004;
ROM_DATA[14] = 32'hafa30008;
ROM_DATA[15] = 32'hafa4000c;
ROM_DATA[16] = 32'hafa50010;
ROM_DATA[17] = 32'hafa60014;
ROM_DATA[18] = 32'hafa70018;
ROM_DATA[19] = 32'hafa8001c;
ROM_DATA[20] = 32'hafa90020;
ROM_DATA[21] = 32'hafaa0024;
ROM_DATA[22] = 32'hafab0028;
ROM_DATA[23] = 32'hafac002c;
ROM_DATA[24] = 32'hafad0030;
ROM_DATA[25] = 32'hafae0034;
ROM_DATA[26] = 32'hafaf0038;
ROM_DATA[27] = 32'hafb0003c;
ROM_DATA[28] = 32'hafb10040;
ROM_DATA[29] = 32'hafb20044;
ROM_DATA[30] = 32'hafb30048;
ROM_DATA[31] = 32'hafb4004c;
ROM_DATA[32] = 32'hafb50050;
ROM_DATA[33] = 32'hafb60054;
ROM_DATA[34] = 32'hafb70058;
ROM_DATA[35] = 32'hafb8005c;
ROM_DATA[36] = 32'hafb90060;
ROM_DATA[37] = 32'hafba0064;
ROM_DATA[38] = 32'hafbb0068;
ROM_DATA[39] = 32'hafbc006c;
ROM_DATA[40] = 32'hafbd0070;
ROM_DATA[41] = 32'hafbe0074;
ROM_DATA[42] = 32'hafbf0078;
ROM_DATA[43] = 32'h27bd007c;
ROM_DATA[44] = 32'h0c000092;
ROM_DATA[45] = 32'h27bdff84;
ROM_DATA[46] = 32'h8fa10000;
ROM_DATA[47] = 32'h8fa20004;
ROM_DATA[48] = 32'h8fa30008;
ROM_DATA[49] = 32'h8fa4000c;
ROM_DATA[50] = 32'h8fa50010;
ROM_DATA[51] = 32'h8fa60014;
ROM_DATA[52] = 32'h8fa70018;
ROM_DATA[53] = 32'h8fa8001c;
ROM_DATA[54] = 32'h8fa90020;
ROM_DATA[55] = 32'h8faa0024;
ROM_DATA[56] = 32'h8fab0028;
ROM_DATA[57] = 32'h8fac002c;
ROM_DATA[58] = 32'h8fad0030;
ROM_DATA[59] = 32'h8fae0034;
ROM_DATA[60] = 32'h8faf0038;
ROM_DATA[61] = 32'h8fb0003c;
ROM_DATA[62] = 32'h8fb10040;
ROM_DATA[63] = 32'h8fb20044;
ROM_DATA[64] = 32'h8fb30048;
ROM_DATA[65] = 32'h8fb4004c;
ROM_DATA[66] = 32'h8fb50050;
ROM_DATA[67] = 32'h8fb60054;
ROM_DATA[68] = 32'h8fb70058;
ROM_DATA[69] = 32'h8fb8005c;
ROM_DATA[70] = 32'h8fb90060;
ROM_DATA[71] = 32'h8fba0064;
ROM_DATA[72] = 32'h8fbb0068;
ROM_DATA[73] = 32'h8fbc006c;
ROM_DATA[74] = 32'h8fbd0070;
ROM_DATA[75] = 32'h8fbe0074;
ROM_DATA[76] = 32'h8fbf0078;
ROM_DATA[77] = 32'h275afffc;
ROM_DATA[78] = 32'h03400008;
ROM_DATA[79] = 32'hafa10000;
ROM_DATA[80] = 32'hafa20004;
ROM_DATA[81] = 32'hafa30008;
ROM_DATA[82] = 32'hafa4000c;
ROM_DATA[83] = 32'hafa50010;
ROM_DATA[84] = 32'hafa60014;
ROM_DATA[85] = 32'hafa70018;
ROM_DATA[86] = 32'hafa8001c;
ROM_DATA[87] = 32'hafa90020;
ROM_DATA[88] = 32'hafaa0024;
ROM_DATA[89] = 32'hafab0028;
ROM_DATA[90] = 32'hafac002c;
ROM_DATA[91] = 32'hafad0030;
ROM_DATA[92] = 32'hafae0034;
ROM_DATA[93] = 32'hafaf0038;
ROM_DATA[94] = 32'hafb0003c;
ROM_DATA[95] = 32'hafb10040;
ROM_DATA[96] = 32'hafb20044;
ROM_DATA[97] = 32'hafb30048;
ROM_DATA[98] = 32'hafb4004c;
ROM_DATA[99] = 32'hafb50050;
ROM_DATA[100] = 32'hafb60054;
ROM_DATA[101] = 32'hafb70058;
ROM_DATA[102] = 32'hafb8005c;
ROM_DATA[103] = 32'hafb90060;
ROM_DATA[104] = 32'hafba0064;
ROM_DATA[105] = 32'hafbb0068;
ROM_DATA[106] = 32'hafbc006c;
ROM_DATA[107] = 32'hafbd0070;
ROM_DATA[108] = 32'hafbe0074;
ROM_DATA[109] = 32'hafbf0078;
ROM_DATA[110] = 32'h27bd007c;
ROM_DATA[111] = 32'h0c000097;
ROM_DATA[112] = 32'h27bdff84;
ROM_DATA[113] = 32'h8fa10000;
ROM_DATA[114] = 32'h8fa20004;
ROM_DATA[115] = 32'h8fa30008;
ROM_DATA[116] = 32'h8fa4000c;
ROM_DATA[117] = 32'h8fa50010;
ROM_DATA[118] = 32'h8fa60014;
ROM_DATA[119] = 32'h8fa70018;
ROM_DATA[120] = 32'h8fa8001c;
ROM_DATA[121] = 32'h8fa90020;
ROM_DATA[122] = 32'h8faa0024;
ROM_DATA[123] = 32'h8fab0028;
ROM_DATA[124] = 32'h8fac002c;
ROM_DATA[125] = 32'h8fad0030;
ROM_DATA[126] = 32'h8fae0034;
ROM_DATA[127] = 32'h8faf0038;
ROM_DATA[128] = 32'h8fb0003c;
ROM_DATA[129] = 32'h8fb10040;
ROM_DATA[130] = 32'h8fb20044;
ROM_DATA[131] = 32'h8fb30048;
ROM_DATA[132] = 32'h8fb4004c;
ROM_DATA[133] = 32'h8fb50050;
ROM_DATA[134] = 32'h8fb60054;
ROM_DATA[135] = 32'h8fb70058;
ROM_DATA[136] = 32'h8fb8005c;
ROM_DATA[137] = 32'h8fb90060;
ROM_DATA[138] = 32'h8fba0064;
ROM_DATA[139] = 32'h8fbb0068;
ROM_DATA[140] = 32'h8fbc006c;
ROM_DATA[141] = 32'h8fbd0070;
ROM_DATA[142] = 32'h8fbe0074;
ROM_DATA[143] = 32'h8fbf0078;
ROM_DATA[144] = 32'h275afffc;
ROM_DATA[145] = 32'h03400008;
ROM_DATA[146] = 32'h27a8ff84;
ROM_DATA[147] = 32'h8d1b0068;
ROM_DATA[148] = 32'h33680001;
ROM_DATA[149] = 32'h10080007;
ROM_DATA[150] = 32'h080000e3;
ROM_DATA[151] = 32'h3c084000;
ROM_DATA[152] = 32'h8d080010;
ROM_DATA[153] = 32'h31080002;
ROM_DATA[154] = 32'h14080001;
ROM_DATA[155] = 32'h08000097;
ROM_DATA[156] = 32'h03e00008;
ROM_DATA[157] = 32'h3c08ffff;
ROM_DATA[158] = 32'h3508fff9;
ROM_DATA[159] = 32'h3c094000;
ROM_DATA[160] = 32'h8d2a0008;
ROM_DATA[161] = 32'h01485024;
ROM_DATA[162] = 32'had2a0008;
ROM_DATA[163] = 32'h2409003f;
ROM_DATA[164] = 32'hafa90000;
ROM_DATA[165] = 32'h24090006;
ROM_DATA[166] = 32'hafa90004;
ROM_DATA[167] = 32'h2409005b;
ROM_DATA[168] = 32'hafa90008;
ROM_DATA[169] = 32'h2409004f;
ROM_DATA[170] = 32'hafa9000c;
ROM_DATA[171] = 32'h24090066;
ROM_DATA[172] = 32'hafa90010;
ROM_DATA[173] = 32'h2409006d;
ROM_DATA[174] = 32'hafa90014;
ROM_DATA[175] = 32'h2409007d;
ROM_DATA[176] = 32'hafa90018;
ROM_DATA[177] = 32'h24090007;
ROM_DATA[178] = 32'hafa9001c;
ROM_DATA[179] = 32'h2409007f;
ROM_DATA[180] = 32'hafa90020;
ROM_DATA[181] = 32'h2409006f;
ROM_DATA[182] = 32'hafa90024;
ROM_DATA[183] = 32'h2409006f;
ROM_DATA[184] = 32'hafa90028;
ROM_DATA[185] = 32'h2409007c;
ROM_DATA[186] = 32'hafa9002c;
ROM_DATA[187] = 32'h24090039;
ROM_DATA[188] = 32'hafa90030;
ROM_DATA[189] = 32'h2409005e;
ROM_DATA[190] = 32'hafa90034;
ROM_DATA[191] = 32'h2409007b;
ROM_DATA[192] = 32'hafa90038;
ROM_DATA[193] = 32'h24090071;
ROM_DATA[194] = 32'hafa9003c;
ROM_DATA[195] = 32'h3c124000;
ROM_DATA[196] = 32'h8e4a0014;
ROM_DATA[197] = 32'h31480f00;
ROM_DATA[198] = 32'h00088242;
ROM_DATA[199] = 32'h14100001;
ROM_DATA[200] = 32'h24100008;
ROM_DATA[201] = 32'h240a0001;
ROM_DATA[202] = 32'h240b0002;
ROM_DATA[203] = 32'h240c0004;
ROM_DATA[204] = 32'h1150000a;
ROM_DATA[205] = 32'h11700006;
ROM_DATA[206] = 32'h11900003;
ROM_DATA[207] = 32'h309100f0;
ROM_DATA[208] = 32'h00118902;
ROM_DATA[209] = 32'h080000d8;
ROM_DATA[210] = 32'h3091000f;
ROM_DATA[211] = 32'h080000d8;
ROM_DATA[212] = 32'h30b100f0;
ROM_DATA[213] = 32'h00118902;
ROM_DATA[214] = 32'h080000d8;
ROM_DATA[215] = 32'h30b1000f;
ROM_DATA[216] = 32'h00115080;
ROM_DATA[217] = 32'h03aa5020;
ROM_DATA[218] = 32'h8d4a0000;
ROM_DATA[219] = 32'h00104200;
ROM_DATA[220] = 32'h010a1020;
ROM_DATA[221] = 32'hae420014;
ROM_DATA[222] = 32'h3c094000;
ROM_DATA[223] = 32'h8d2a0008;
ROM_DATA[224] = 32'h354a0002;
ROM_DATA[225] = 32'had2a0008;
ROM_DATA[226] = 32'h0800009c;
ROM_DATA[227] = 32'h3c104000;
ROM_DATA[228] = 32'h8e090020;
ROM_DATA[229] = 32'h31290004;
ROM_DATA[230] = 32'h1009fffc;
ROM_DATA[231] = 32'h8e080018;
ROM_DATA[232] = 32'h0800009c;

end
endmodule
